library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity TheirVGA is
port(mclk: in std_logic;
        ledvga: in std_logic_vector(14 downto 0);
        modev: in std_logic;
        modev2: in std_logic;
        TLv: in std_logic_vector(15 downto 0);
        TSv: in std_logic_vector(15 downto 0);
        timeremain1: in std_logic_vector(15 downto 0);
		vs, hs: out std_logic;
		red, grn, blu : out std_logic_vector(3 downto 0));
end TheirVGA;

architecture Behavioral of TheirVGA is
signal clkPix: std_logic;
signal cntHorz, cntVert: std_logic_vector(9 downto 0);
signal charpixcount1, charpixcount2: integer:=0;
signal sncHorz, clkLine, blkHorz, sncVert, blkVert, blkDisp, clkColor: std_logic;
signal cntImg: std_logic_vector(6 downto 0);
--signal cntColor: std_logic_vector(11 downto 0);
signal cntColor: std_logic_vector(11 downto 0);
signal cntColor1: std_logic_vector(11 downto 0);
signal nrcolor,nycolor,ngcolor,nacolor,srcolor,sycolor,sgcolor,sacolor,ercolor,eycolor,egcolor,eacolor,wrcolor,wycolor,wgcolor,wacolor: std_logic_vector(11 downto 0);
signal sercolor,seycolor,segcolor:std_logic_vector(11 downto 0); 
signal upper, left, lower, right: std_logic_vector(11 downto 0);
signal tnr,tny,tng,tna,tsr,tsy,tsg,tsa,ter,tey,teg,tea,twr,twy,twg,twa,tser,tsey,tseg: std_logic_vector(11 downto 0);
signal bnr,bny,bng,bna,bsr,bsy,bsg,bsa,ber,bey,beg,bea,bwr,bwy,bwg,bwa,bser,bsey,bseg: std_logic_vector(11 downto 0);
signal lnr,lny,lng,lna,lsr,lsy,lsg,lsa,ler,ley,leg,lea,lwr,lwy,lwg,lwa,lser,lsey,lseg: std_logic_vector(11 downto 0);
signal rnr,rny,rng,rna,rsr,rsy,rsg,rsa,rer,rey,reg,rea,rwr,rwy,rwg,rwa,rser,rsey,rseg: std_logic_vector(11 downto 0);
signal tsec0,bsec0,lsec0,rsec0,tsec1,bsec1,lsec1,rsec1:std_logic_vector(11 downto 0);
signal count: std_logic_vector(1 downto 0);
type char_type is array (0 to 31) of std_logic_vector(0 to 31); --32x32 character resolution
signal value0: char_type;
signal value1: char_type;

constant zero: char_type:= (
"00000000000011111111100000000000",
"00000000001111111111111000000000",
"00000000111111111111111110000000",
"00000001111111111111111111000000",
"00000011111111111111111111100000",
"00000111111111000001111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111110000000111111110000",
"00000111111111000001111111110000",
"00000011111111111111111111100000",
"00000001111111111111111111000000",
"00000000111111111111111110000000",
"00000000001111111111111000000000",
"00000000000011111111100000000000"
);

constant one: char_type:= (
"00000000000011111111000000000000",
"00000000000111111111000000000000",
"00000000001111111111000000000000",
"00000000011111111111000000000000",
"00000000111111111111000000000000",
"00000001111111111111000000000000",
"00000011111111111111000000000000",
"00000111111111111111000000000000",
"00001111111111111111000000000000",
"00001111111111111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00001111111111111111111111110000"
);

constant two: char_type:= (
"00000000000011111111000000000000",
"00000000001111111111110000000000",
"00000000111111111111111100000000",
"00000011111111111111111111000000",
"00000111111111111111111111100000",
"00001111111111111111111111110000",
"00011111111111111111111111111000",
"00011111111110000000111111111100",
"00111111111100000000011111111100",
"00111111111000000000011111111110",
"01111111110000000000011111111110",
"01111111110000000000011111111110",
"01111111110000000000111111111110",
"00000000000000000001111111111110",
"00000000000000000011111111111110",
"00000000000000000111111111111100",
"00000000000000011111111111111100",
"00000000000001111111111111111000",
"00000000000011111111111111110000",
"00000000001111111111111111100000",
"00000000111111111111111111000000",
"00000001111111111111111110000000",
"00000111111111111111111000000000",
"00001111111111111111110000000000",
"00011111111111111111000000000000",
"00111111111111111100000000000000",
"00111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110"
);

constant three: char_type:= (
"00000000000011111111111100000000",
"00000000001111111111111111000000",
"00000000111111111111111111100000",
"00000011111111111111111111110000",
"00000111111111111111111111111000",
"00001111111111111111111111111100",
"00011111111111111111111111111100",
"00011111111110000000111111111110",
"00111111111100000000011111111110",
"00111111111000000000011111111110",
"01111111110000000000011111111110",
"00000000000000000000011111111110",
"00000000000000000000111111111110",
"00000000000000011111111111111100",
"00000000000000011111111111111000",
"00000000000000011111111111100000",
"00000000000000011111111111111000",
"00000000000000011111111111111100",
"00000000000000011111111111111110",
"00000000000000000000111111111110",
"00000000000000000000011111111110",
"01111111110000000000011111111110",
"00111111111000000000011111111110",
"00111111111100000000011111111110",
"00011111111110000000111111111100",
"00011111111111111111111111111100",
"00001111111111111111111111111000",
"00000111111111111111111111110000",
"00000011111111111111111111100000",
"00000001111111111111111111000000",
"00000000011111111111111110000000",
"00000000000111111111111000000000"
);

constant four: char_type:= (
"00000000000000000011111111110000",
"00000000000000000111111111110000",
"00000000000000001111111111110000",
"00000000000000011111111111110000",
"00000000000000111111111111110000",
"00000000000001111111111111110000",
"00000000000011111111111111110000",
"00000000000111111111111111110000",
"00000000001111111111111111110000",
"00000000011111111101111111110000",
"00000000111111111001111111110000",
"00000001111111110001111111110000",
"00000011111111100001111111110000",
"00000111111111000001111111110000",
"00001111111110000001111111110000",
"00011111111100000001111111110000",
"00111111111000000001111111110000",
"01111111110000000001111111110000",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"00000000000000000001111111110000",
"00000000000000000001111111110000",
"00000000000000000001111111110000",
"00000000000000000001111111110000",
"00000000000000000001111111110000"
);

constant five: char_type:= (
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111000000000001111111110",
"01111111111000000000001111111110",
"01111111111000000000001111111110",
"01111111111000000000001111111110",
"01111111111000000000000000000000",
"01111111111000000000000000000000",
"01111111111111111111111111000000",
"01111111111111111111111111110000",
"01111111111111111111111111111000",
"01111111111111111111111111111100",
"01111111111111111111111111111100",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"00000000000000000000111111111110",
"00000000000000000000011111111110",
"00000000000000000000011111111110",
"00000000000000000000011111111110",
"01111111111100000000011111111110",
"01111111111110000000111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"00111111111111111111111111111100",
"00111111111111111111111111111100",
"00011111111111111111111111111000",
"00001111111111111111111111110000",
"00000011111111111111111111000000"
);

constant six: char_type:= (
"00000011111111111111111111000000",
"00001111111111111111111111110000",
"00011111111111111111111111111000",
"00111111111111111111111111111100",
"00111111111111111111111111111100",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111110000000111111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111100000000000000000000",
"01111111111100000000000000000000",
"01111111111110000000000000000000",
"01111111111111111111111111100000",
"01111111111111111111111111111000",
"01111111111111111111111111111100",
"01111111111111111111111111111100",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111110000000111111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111110000000111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"00111111111111111111111111111100",
"00111111111111111111111111111100",
"00011111111111111111111111111000",
"00001111111111111111111111110000",
"00000011111111111111111111000000"
);

constant seven: char_type:= (
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111110000000000001111111110",
"01111111110000000000001111111110",
"01111111110000000000001111111110",
"00000000000000000000001111111110",
"00000000000000000000011111111100",
"00000000000000000000111111111000",
"00000000000000000001111111110000",
"00000000000000000011111111100000",
"00000000000000000111111111000000",
"00000000000000001111111110000000",
"00000000000000011111111100000000",
"00000000000000111111111000000000",
"00000000000001111111110000000000",
"00000000000011111111100000000000",
"00000000000111111111000000000000",
"00000000001111111110000000000000",
"00000000011111111100000000000000",
"00000000111111111000000000000000",
"00000001111111110000000000000000",
"00000011111111100000000000000000",
"00000111111111000000000000000000",
"00001111111110000000000000000000",
"00011111111100000000000000000000",
"00111111111000000000000000000000",
"01111111110000000000000000000000",
"01111111110000000000000000000000"
);

constant eight: char_type:= (
"00000011111111111111111111000000",
"00001111111111111111111111110000",
"00011111111111111111111111111000",
"00111111111111111111111111111100",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111110000000111111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111110000000111111111110",
"00111111111111111111111111111100",
"00011111111111111111111111111000",
"00000111111111111111111111100000",
"00011111111111111111111111111000",
"00111111111111111111111111111100",
"01111111111111111111111111111110",
"01111111111110000000111111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111110000000111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"00111111111111111111111111111100",
"00111111111111111111111111111100",
"00011111111111111111111111111000",
"00001111111111111111111111110000",
"00000011111111111111111111000000"

);

constant nine: char_type:= (
"00000011111111111111111111000000",
"00001111111111111111111111110000",
"00011111111111111111111111111000",
"00111111111111111111111111111100",
"00111111111111111111111111111100",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111110000000111111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111100000000011111111110",
"01111111111110000000111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"00111111111111111111111111111110",
"00111111111111111111111111111110",
"00011111111111111111111111111110",
"00000111111111111111111111111110",
"00000000000000000000111111111110",
"00000000000000000000011111111110",
"00000000000000000000011111111110",
"00000000000000000000011111111110",
"01111111111100000000011111111110",
"01111111111110000000111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"00111111111111111111111111111100",
"00111111111111111111111111111100",
"00011111111111111111111111111000",
"00001111111111111111111111110000",
"00000011111111111111111111000000"
);

constant light: char_type:= (
"00000000000011111111000000000000",
"00000000001111111111110000000000",
"00000000111111111111111100000000",
"00000011111111111111111111000000",
"00000111111111111111111111100000",
"00001111111111111111111111110000",
"00011111111111111111111111111000",
"00011111111111111111111111111000",
"00111111111111111111111111111100",
"00111111111111111111111111111100",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"11111111111111111111111111111111",
"11111111111111111111111111111111",
"11111111111111111111111111111111",
"11111111111111111111111111111111",
"11111111111111111111111111111111",
"11111111111111111111111111111111",
"11111111111111111111111111111111",
"11111111111111111111111111111111",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"00111111111111111111111111111100",
"00111111111111111111111111111100",
"00011111111111111111111111111000",
"00011111111111111111111111111000",
"00001111111111111111111111110000",
"00000111111111111111111111100000",
"00000011111111111111111111000000",
"00000000111111111111111100000000",
"00000000001111111111110000000000",
"00000000000011111111000000000000"
);

constant na: char_type:= (
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"11111111111111000000000000000000",
"11111111111111000000000000000000",
"11111111111111000000000000000000",
"11111111111111000000000000000000",
"11111111111111000000000000000000",
"11111111111111000000000000000000",
"11111111111111000000000000000000",
"11111111111111000000000000000000",
"11111111111111000000000000000000",
"11111111111111000000000000000000",
"11111111111111000000000100000000",
"11111111111111000000000110000000",
"11111111111111000000000111000000",
"11111111111111000000000111100000",
"11111111111111111111111111110000",
"11111111111111111111111111111000",
"11111111111111111111111111111100",
"11111111111111111111111111111110",
"11111111111111111111111111111111",
"11111111111111111111111111111110",
"11111111111111111111111111111100",
"11111111111111111111111111111000",
"11111111111111111111111111110000",
"00000000000000000000000111100000",
"00000000000000000000000111000000",
"00000000000000000000000110000000",
"00000000000000000000000100000000",
"00000000000000000000000000000000"
);

constant sa: char_type:= (
"00000000010000000000000000000000",
"00000000110000000000000000000000",
"00000001110000000000000000000000",
"00000011110000000000000000000000",
"00000111110000000000000000000000",
"00001111111111111111111111111111",
"00011111111111111111111111111111",
"00111111111111111111111111111111",
"01111111111111111111111111111111",
"11111111111111111111111111111111",
"01111111111111111111111111111111",
"00111111111111111111111111111111",
"00011111111111111111111111111111",
"00001111111111111111111111111111",
"00000111110000000001111111111111",
"00000011110000000000111111111111",
"00000001110000000000011111111111",
"00000000110000000000001111111111",
"00000000010000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111",
"00000000000000000000000111111111"
);

constant wa: char_type:= (
"00000000000000000000001000000000",
"00000000000000000000011100000000",
"00000000000000000000111110000000",
"00000000000000000001111111000000",
"00000000000000000011111111100000",
"00000000000000000111111111110000",
"00000000000000001111111111111000",
"00000000000000011111111111111100",
"00000000000000111111111111111110",
"00000000000001111111111111111111",
"00000000000000000011111111100000",
"00000000000000000011111111100000",
"00000000000000000011111111100000",
"00000000000000000011111111100000",
"00000000000000000011111111100000",
"00000000000000000011111111100000",
"00000000000000000011111111100000",
"00000000000000000011111111100000",
"00000000000000000011111111100000",
"00000000000000000111111111100000",
"00000000000000001111111111100000",
"00000000000000011111111111100000",
"00000000000000111111111111100000",
"11111111111111111111111111100000",
"11111111111111111111111111100000",
"11111111111111111111111111100000",
"11111111111111111111111111100000",
"11111111111111111111111111100000",
"11111111111111111111111111100000",
"11111111111111111111111111100000",
"11111111111111111111111111100000",
"11111111111111111111111111100000"
);

constant ea: char_type:= (
"00000111111111111111111111111111",
"00000111111111111111111111111111",
"00000111111111111111111111111111",
"00000111111111111111111111111111",
"00000111111111111111111111111111",
"00000111111111111111111111111111",
"00000111111111111111111111111111",
"00000111111111111111111111111111",
"00000111111111111111111111111111",
"00000111111111111100000000000000",
"00000111111111111000000000000000",
"00000111111111110000000000000000",
"00000111111111100000000000000000",
"00000111111111000000000000000000",
"00000111111111000000000000000000",
"00000111111111000000000000000000",
"00000111111111000000000000000000",
"00000111111111000000000000000000",
"00000111111111000000000000000000",
"00000111111111000000000000000000",
"00000111111111000000000000000000",
"00000111111111000000000000000000",
"11111111111111111110000000000000",
"01111111111111111100000000000000",
"00111111111111111000000000000000",
"00011111111111110000000000000000",
"00001111111111100000000000000000",
"00000111111111000000000000000000",
"00000011111110000000000000000000",
"00000001111100000000000000000000",
"00000000111000000000000000000000",
"00000000010000000000000000000000"
);

constant tee: char_type:= (
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000",
"00000000000011111111000000000000");

constant el: char_type:= (
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111100000000000000000000000",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110");

constant ess: char_type:= (
"00000011111111111111111111000000",
"00001111111111111111111111110000",
"00011111111111111111111111111000",
"00111111111111111111111111111100",
"00111111111111111111111111111100",
"01111111111111111111111111111110",
"01111111111100000000011111111110",
"01111111111000000000001111111110",
"01111111111000000000001111111110",
"01111111111000000000001111111110",
"01111111111000000000000000000000",
"01111111111100000000000000000000",
"01111111111111111111111111000000",
"01111111111111111111111111110000",
"00111111111111111111111111111000",
"00111111111111111111111111111100",
"00011111111111111111111111111100",
"00001111111111111111111111111110",
"00000011111111111111111111111110",
"00000000000000000000111111111110",
"00000000000000000000011111111110",
"00000000000000000000011111111110",
"00000000000000000000011111111110",
"01111111111100000000011111111110",
"01111111111110000000111111111110",
"01111111111111111111111111111110",
"01111111111111111111111111111110",
"00111111111111111111111111111100",
"00111111111111111111111111111100",
"00011111111111111111111111111000",
"00001111111111111111111111110000",
"00000011111111111111111111000000");

constant equal: char_type:= (
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00001111111111111111111111110000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000");


begin

tnr<=X"01B"; --north red
bnr<=X"03B";
lnr<=X"19A";
rnr<=X"1BA";

tny<=bnr+3; --north yellow
bny<=tny+32;
lny<=X"19A";
rny<=X"1BA";

tng<=bny+3; --north green
bng<=tng+32;
lng<=X"19A";
rng<=X"1BA";

tna<=tng; --north arrow
bna<=bng;
lna<=rng+3;
rna<=lna+32;

tsr<=tng+350; --south red
bsr<=bng+350;
lsr<=X"19A";
rsr<=X"1BA";

tsy<=tny+350; --south yellow
bsy<=bny+350;
lsy<=X"19A";
rsy<=X"1BA";

tsg<=tnr+350; --south green
bsg<=bnr+350;
lsg<=X"19A";
rsg<=X"1BA";

tsa<=tsg; --south arrow
bsa<=bsg;
lsa<=lsg-35;
rsa<=lsa+32;

twr<=X"0D8"; --west red
bwr<=twr+32;
lwr<=X"0A5";
rwr<=lwr+32;

twy<=twr; --west yellow
bwy<=bwr;
lwy<=rwr+3;
rwy<=lwy+32;

twg<=twr; --west green
bwg<=bwr;
lwg<=rwy+3;
rwg<=lwg+32;

twa<=twg-35; --west arrow
bwa<=twa+32;
lwa<=lwg;
rwa<=rwg;

ter<=twr; --east red
ber<=bwr;
ler<=lwg+430;
rer<=ler+32;

tey<=twr; --east yellow
bey<=bwr;
ley<=lwy+430;
rey<=ley+32;

teg<=twr; --east green
beg<=bwr;
leg<=lwr+430;
reg<=leg+32;

tea<=teg+35; --east arrow
bea<=tea+32;
lea<=leg;
rea<=reg;

tsec1<=teg; --left secs digit
bsec1<=beg;
lsec1<=lng;
rsec1<=rng;

tsec0<=teg; --right secs digit
bsec0<=beg;
lsec0<=lna;
rsec0<=rna;

tser<=tsr; --southeast red
bser<=bsr;
lser<=ler;
rser<=rer;

tsey<=tsy; --southeast yellow
bsey<=bsy;
lsey<=ley;
rsey<=rey;

tseg<=tsg; --southeast green
bseg<=bsg;
lseg<=leg;
rseg<=reg;

------------------------------------------------------------------------
    --          VGA Controller Test
	------------------------------------------------------------------------

    -- Divide the D2XL oscillator down to form the pixel clock
    -- that is the basis for all of the other timing.
    process (mclk)
        begin
            if mclk = '1' and mclk'Event then
            if (count = "10") then
                count <= "00";
                clkPix <= not clkPix;
            else
                count <= count+1;
            end if;
            end if;
        end process;

    -- Generate the horizontal timing.
    process (clkPix)
        begin
		  		
            if clkPix = '1' and clkPix'Event then
                if cntHorz = "0001011101" then  -- horizontal sync pulse is 93 pixels long
                    cntHorz <= cntHorz + 1; --increment pixel count
                    sncHorz <= '1'; -- back porch starts here, turn on horizontal sync signal
                elsif cntHorz = "0010001100" then --140: start of video display section (after horizontal sync pulse and back porch)
                    cntHorz <= cntHorz + 1; 
                    blkHorz <= '0'; --video on
                elsif cntHorz = "1100001100" then --780: end of video display section(780-140=640 pixels) 
                    cntHorz <= cntHorz + 1;
                    blkHorz <= '1'; --video off
                elsif cntHorz = "1100011010" then --794: end of horizontal line (14 pixels for front porch)
                    cntHorz <= "0000000000"; --reset horizontal pixel count
                    clkLine <= '1'; -- set clock signal for vertical timing
                    sncHorz <= '0'; -- pulse horizontal sync low to indicate beginning of next horizontal line
                else
                    cntHorz <= cntHorz + 1;
                    clkLine <= '0';
                end if;
            end if;
        end process;

    -- Generate the vertical timing.
    process (clkLine)
        begin
		  		
            if clkLine = '1' and clkLine'Event then
                if cntVert = "0000000001" then --vertical sync pulse is 2 pixel long
                    cntVert <= cntVert + 1; --increment line/row count by 1
                    sncVert <= '1'; -- vertical back porch starts here, sent vertical sync signal high
                elsif cntVert = "0000011010" then --26: end of vertical back porch; beginning of video display section
                    cntVert <= cntVert + 1;
                    blkVert <= '0'; --video on
                elsif cntVert = "0111111010" then --506: end of video display section
                    cntVert <= cntVert + 1;
                    blkVert <= '1'; --video off
                elsif cntVert = "1000001100" then -- 524: end of frame (front porch is 18 pixels long)
                    cntVert <= "0000000000"; -- reset line/row count
                    sncVert <= '0'; -- pulse vertical sync signal to indicate beginning of new frame
                   else
               
                cntVert <= cntVert + 1; --increment line/row count
          end if;
          end if;
          
        end process;
        
        process(clkpix)
        begin
          if clkPix = '1' and clkPix'Event then
            if (cntHorz>lnr and cntHorz<rnr)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lny and cntHorz<rny)then
             charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lng and cntHorz<rng)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lna and cntHorz<rna)then
            charpixcount1<=charpixcount1+1;
            elsif(cntHorz>lsr and cntHorz<rsr)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lsy and cntHorz<rsy)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lsg and cntHorz<rsg)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lsa and cntHorz<rsa)then
            charpixcount1<=charpixcount1+1;
            elsif(cntHorz>ler and cntHorz<rer)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>ley and cntHorz<rey)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>leg and cntHorz<reg)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lea and cntHorz<rea)then
            charpixcount1<=charpixcount1+1;
            elsif(cntHorz>lwr and cntHorz<rwr)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lwy and cntHorz<rwy)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lwg and cntHorz<rwg)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lwa and cntHorz<rwa)then
            charpixcount1<=charpixcount1+1;
            elsif(cntHorz>lser and cntHorz<rser)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lsey and cntHorz<rsey)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lseg and cntHorz<rseg)then
            charpixcount1<=charpixcount1+1;
             elsif(cntHorz>lsec0 and cntHorz<rsec0)then
             charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lsec1 and cntHorz<rsec1)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lsec1-70 and cntHorz<rsec1-70)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lsec1-35 and cntHorz<rsec1-35)then
            charpixcount1<=charpixcount1+1;
            elsif (cntHorz>lsec1+70 and cntHorz<rsec1+70)then
            charpixcount1<=charpixcount1+1;
            else
            charpixcount1<=0;
            end if;
        end if;
        end process;
        
         process(clkLine)
               begin
                 if clkLine = '1' and clkLine'Event then
                   if (cntVert>tnr and cntVert<bnr)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tny and cntVert<bny)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tng and cntVert<bng)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tna and cntVert<bna)then
                   charpixcount2<=charpixcount2+1;
                   elsif(cntVert>tsr and cntVert<bsr)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tsy and cntVert<bsy)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tsg and cntVert<bsg)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tsa and cntVert<bsa)then
                   charpixcount2<=charpixcount2+1;
                   elsif(cntVert>ter and cntVert<ber)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tey and cntVert<bey)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>teg and cntVert<beg)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tea and cntVert<bea)then
                   charpixcount2<=charpixcount2+1;
                   elsif(cntVert>twr and cntVert<bwr)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>twy and cntVert<bwy)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>twg and cntVert<bwg)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>twa and cntVert<bwa)then
                   charpixcount2<=charpixcount2+1;
                   elsif(cntVert>tser and cntVert<bser)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tsey and cntVert<bsey)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tseg and cntVert<bseg) then
                   charpixcount2<=charpixcount2+1;
                   elsif(cntVert>tsec0 and cntVert<bsec0)then
                   charpixcount2<=charpixcount2+1;
                   elsif (cntVert>tsec1 and cntVert<bsec1)then
                   charpixcount2<=charpixcount2+1;
                   else
                   charpixcount2<=0;
                   end if;
               end if;
               end process;
               
               process(timeremain1)
               begin
             if(mclk'event and mclk='1') then
             if modev='0' then
               if timeremain1="0010011100010000" then   --10000 for 10secs
                value0<=zero;
                value1<=one;
               elsif timeremain1="0010001100101000" then   --9000 for 9secs
                  value0<=nine;
                  value1<=zero;
              elsif timeremain1="0001111101000000" then   --8000 for 8secs
                 value0<=eight;
                 value1<=zero;
              elsif timeremain1="0001101101011000" then   --7000 for 7secs
                value0<=seven;
                value1<=zero;
               elsif timeremain1="0001011101110000" then   --6000 for 6secs
                value0<=six;
                value1<=zero;
               elsif timeremain1="0001001110001000" then   --5000 for 5secs
                   value0<=five;
                   value1<=zero;
               elsif timeremain1="0000111110100000" then   --4000 for 4secs
                    value0<=four;
                    value1<=zero;
                elsif timeremain1="0000101110111000" then   --3000 for 3secs
                    value0<=three;
                    value1<=zero;
                elsif timeremain1="0000011111010000" then   --2000 for 2secs
                    value0<=two;
                    value1<=zero;
                elsif timeremain1="0000001111101000" then   --1000 for 1sec
                   value0<=one;
                   value1<=zero;
                elsif timeremain1="0000000000000000" then   --0 for 0secs
                   value0<=zero;
                   value1<=zero;
                end if;
             else
                if modev2='0' then
                           if TLv="0010011100010000" then   --10secs
                             value0<=zero;
                             value1<=one;
                            elsif TLv="0010001100101000" then   --9secs
                               value0<=nine;
                               value1<=zero;
                           elsif TLv="0001111101000000" then   --8secs
                              value0<=eight;
                              value1<=zero;
                           elsif TLv="0001101101011000" then   --7secs
                             value0<=seven;
                             value1<=zero;
                            elsif TLv="0001011101110000"  then   --6secs
                             value0<=six;
                             value1<=zero;
                            elsif TLv="0001001110001000" then   --5secs
                                value0<=five;
                                value1<=zero;
                            elsif TLv="0000111110100000" then   --4secs
                                 value0<=four;
                                 value1<=zero;
                             elsif TLv="0000101110111000" then   -- 3secs
                                 value0<=three;
                                 value1<=zero;
                             elsif TLv="0000011111010000" then   -- 2secs
                                 value0<=two;
                                 value1<=zero;
                             elsif TLv="0000001111101000" then   -- 1sec
                                value0<=one;
                                value1<=zero;
                             elsif TLv="0000000000000000" then   -- 0secs
                                value0<=zero;
                                value1<=zero;
                           end if;
                         if TSv="0010011100010000" then   --10secs
                                                     value0<=zero;
                                                      value1<=one;
                                                    elsif TSv="0010001100101000" then   --9secs
                                                      value0<=nine;
                                                       value1<=zero;
                                                  elsif TSv="0001111101000000" then   --8secs
                                                      value0<=eight;
                                                      value1<=zero;
                                                   elsif TSv="0001101101011000" then   --7secs
                                                     value0<=seven;
                                                     value1<=zero;
                                                    elsif TSv="0001011101110000"  then   --6secs
                                                     value0<=six;
                                                     value1<=zero;
                                                    elsif TSv="0001001110001000" then   --5secs
                                                         value0<=five;
                                                         value1<=zero;
                                                    elsif TSv="0000111110100000" then   --4secs
                                                         value0<=four;
                                                          value1<=zero;
                                                     elsif TSv="0000101110111000" then   -- 3secs
                                                         value0<=three;
                                                         value1<=zero;
                                                     elsif TSv="0000011111010000" then   -- 2secs
                                                         value0<=two;
                                                         value1<=zero;
                                                     elsif TSv="0000001111101000" then   -- 1sec
                                                        value0<=one;
                                                        value1<=zero;
                                                     elsif TSv="0000000000000000" then   -- 0secs
                                                        value0<=zero;
                                                         value1<=zero;
                                                    end if;
                                                   end if;
--                
             end if;
             end if;
           end process;
               
   -- Divide the active portion of a scan line into 8 regions.
    -- This counts up to 79 and then resets. Each time it
    -- resets, it generates a pulse on clkColor.
    process (clkPix, blkDisp)
        begin
            if clkPix = '1' and clkPix'Event then
                if blkDisp = '1' then -- video off region
                    cntImg <= "0000000";
                else
                    if cntImg = "1001111" then  --79 pulse signal clkColor after every 79 pixels in "video on" region
                        cntImg <= "0000000";
                        clkColor <= '1';
                    else
                        cntImg <= cntImg + 1;
                        clkColor <= '0';
                    end if;
                end if;
            end if;
        end process;
	
    blkDisp <= blkVert or blkHorz;
    
    process(cntHorz,cntVert)
    begin
    
    if modev='0' then --Display mode
    -- all red lights
    if(cntHorz < rnr and cntHorz > lnr and cntVert < bnr and cntVert > tnr and light(charpixcount2)(charpixcount1)='1')then
        if(ledvga ="110000000000000" or ledvga="100000000000000" or ledvga="111111000000000" or ledvga="101111000000000") then
        cntColor <= "010000000000"; --dim red
        else
        cntColor <= "111100000000"; --bright red
        end if;
    elsif (cntHorz < rsr and cntHorz > lsr and cntVert < bsr and cntVert > tsr and light(charpixcount2)(charpixcount1)='1')then
        if(ledvga="111111000000000" or ledvga="101111000000000" or ledvga="000110000000000" or ledvga="000100000000000") then
        cntColor <= "010000000000"; --dim red
        else
        cntColor <= "111100000000"; --bright red
        end if;
    elsif (cntHorz < rer and cntHorz > ler and cntVert < ber and cntVert > ter and light(charpixcount2)(charpixcount1)='1')then
        if(ledvga="000000111111000" or ledvga="000000101101000" or ledvga="000000110000000" or ledvga="000000100000000") then
        cntColor <= "010000000000"; --dim red
        else
        cntColor <= "111100000000"; --bright red
        end if;
    elsif (cntHorz < rwr and cntHorz > lwr and cntVert < bwr and cntVert > twr and light(charpixcount2)(charpixcount1)='1')then
        if(ledvga="000000111111000" or ledvga="000000101101000" or ledvga="000000000110000" or ledvga="000000000100000") then
        cntColor <= "010000000000"; --dim red
        else
        cntColor <= "111100000000"; --bright red
        end if;
     elsif(cntHorz < rser and cntHorz > lser and cntVert < bser and cntVert > tser and light(charpixcount2)(charpixcount1)='1')then
         if(ledvga="000000000000111" or ledvga="000000000000010") then
         cntColor <= "010000000000"; --dim red
         else
         cntColor <= "111100000000"; --bright red
         end if;
    
   --all yellow lights 
    elsif(cntHorz < rny and cntHorz > lny and cntVert < bny and cntVert > tny and light(charpixcount2)(charpixcount1)='1') then
        if(ledvga="101111000000000") then
            cntColor <= "111111110000"; --bright yellow
            else
            cntColor <= "010001000000"; --dim yellow
            end if;
        elsif (cntHorz < rsy and cntHorz > lsy and cntVert < bsy and cntVert > tsy and light(charpixcount2)(charpixcount1)='1')then
            if(ledvga="000100000000000") then
                cntColor <= "111111110000"; --bright yellow
                else
                cntColor <= "010001000000"; --dim yellow
                end if;
        elsif (cntHorz < rey and cntHorz > ley and cntVert < bey and cntVert > tey and light(charpixcount2)(charpixcount1)='1')then
            if(ledvga="000000101101000") then
                 cntColor <= "111111110000"; --bright yellow
                           else
                           cntColor <= "010001000000"; --dim yellow
                           end if;
        elsif (cntHorz < rwy and cntHorz > lwy and cntVert < bwy and cntVert > twy and light(charpixcount2)(charpixcount1)='1')then
            if(ledvga="000000101101000") then
                cntColor <= "111111110000"; --bright yellow
                                       else
                                       cntColor <= "010001000000"; --dim yellow
                                       end if;
       elsif(cntHorz < rsey and cntHorz > lsey and cntVert < bsey and cntVert > tsey and light(charpixcount2)(charpixcount1)='1')then
      
        if(ledvga="000000000000010") then
       cntColor <= "111111110000"; --bright yellow
                                               else
                                               cntColor <= "010001000000"; --dim yellow
                                               end if;
       
       --all green lights 
     elsif(cntHorz < rng and cntHorz > lng and cntVert < bng and cntVert > tng and light(charpixcount2)(charpixcount1)='1') then
        if(ledvga="110000000000000" or ledvga="100000000000000" or ledvga="111111000000000") then
                cntColor <= "000011110000";   --bright green
                else
                cntColor <= "000001000000";     --dim green
                end if;
     elsif(cntHorz < rsg and cntHorz > lsg and cntVert < bsg and cntVert > tsg and light(charpixcount2)(charpixcount1)='1') then
         if(ledvga="111111000000000" or ledvga="101111000000000" or ledvga="000110000000000") then
                    cntColor <= "000011110000";   --bright green
                    else
                    cntColor <= "000001000000";     --dim green
                    end if;
     elsif(cntHorz < reg and cntHorz > leg and cntVert < beg and cntVert > teg and light(charpixcount2)(charpixcount1)='1') then
        if(ledvga="000000111111000" or ledvga="000000110000000" or ledvga="000000100000000") then
                        cntColor <= "000011110000";   --bright green
                        else
                        cntColor <= "000001000000";     --dim green
                        end if;
    elsif(cntHorz < rwg and cntHorz > lwg and cntVert < bwg and cntVert > twg and light(charpixcount2)(charpixcount1)='1') then
       if(ledvga="000000111111000" or ledvga="000000000110000" or ledvga="000000000100000") then
                            cntColor <= "000011110000";   --bright green
                            else
                            cntColor <= "000001000000";     --dim green
                            end if;
    elsif(cntHorz < rseg and cntHorz > lseg and cntVert < bseg and cntVert > tseg and light(charpixcount2)(charpixcount1)='1') then
           if(ledvga="000000000000111") then
           cntColor <= "000011110000";   --bright green
           else
           cntColor <= "000001000000";     --dim green
           end if;
           
     --all arrow lights          
   elsif(cntHorz < rna and cntHorz > lna and cntVert < bna and cntVert > tna and na(charpixcount2)(charpixcount1)='1') then
   if(ledvga="110000000000000") then
             cntColor <= "000011110000";   --bright green
             elsif(ledvga="100000000000000") then
             cntColor <= "111111110000";  --bright yellow
             else
             cntColor <= "001100110011"; -- grey to signify off
             end if;
   elsif(cntHorz < rsa and cntHorz > lsa and cntVert < bsa and cntVert > tsa and sa(charpixcount2)(charpixcount1)='1') then
    if(ledvga="000110000000000") then
               cntColor <= "000011110000";   --bright green
               elsif(ledvga="000100000000000") then
               cntColor <= "111111110000";  --bright yellow
               else
               cntColor <= "001100110011"; -- grey to signify off
               end if;
   elsif(cntHorz < rea and cntHorz > lea and cntVert < bea and cntVert > tea and ea(charpixcount2)(charpixcount1)='1') then
    if(ledvga="000000110000000") then
                 cntColor <= "000011110000";   --bright green
                 elsif(ledvga="000000100000000") then
                 cntColor <= "111111110000";  --bright yellow
                 else
                 cntColor <= "001100110011"; -- grey to signify off
                 end if;
   elsif(cntHorz < rwa and cntHorz > lwa and cntVert < bwa and cntVert > twa and wa(charpixcount2)(charpixcount1)='1') then
         if(ledvga="000000000110000") then
                    cntColor <= "000011110000";   --bright green
                    elsif(ledvga="000000000100000") then
                    cntColor <= "111111110000";  --bright yellow
                    else
                    cntColor <= "001100110011"; -- grey to signify off
                    end if;
  
  --time remaining digits        
elsif((cntHorz < rsec0 and cntHorz > lsec0 and cntVert < bsec0 and cntVert > tsec0 and value0(charpixcount2)(charpixcount1)='1') 
                    or (cntHorz < rsec1 and cntHorz > lsec1 and cntVert < bsec1 and cntVert > tsec1 and value1(charpixcount2)(charpixcount1)='1')
                    ) then
                    cntColor <= "111111111111";   -- white
                    
  else 
        cntColor <= "000000000000";   --black background
       
    end if;
    
 else --display only time in timer change mode
  if modev2='0' then
    if((cntHorz < rsec0+35 and cntHorz > lsec0+35 and cntVert < bsec0 and cntVert > tsec0 and value0(charpixcount2)(charpixcount1)='1') 
                     or (cntHorz < rsec1+35 and cntHorz > lsec1+35 and cntVert < bsec1 and cntVert > tsec1 and value1(charpixcount2)(charpixcount1)='1')
                     or (cntHorz < rsec1 and cntHorz > lsec1 and cntVert < bsec1 and cntVert > tsec1 and equal(charpixcount2)(charpixcount1)='1')
                     or (cntHorz < rsec1-35 and cntHorz > lsec1-35 and cntVert < bsec1 and cntVert > tsec1 and el(charpixcount2)(charpixcount1)='1')
                     or (cntHorz < rsec1-70 and cntHorz > lsec1-70 and cntVert < bsec1 and cntVert > tsec1 and tee(charpixcount2)(charpixcount1)='1')
                     ) then
                     cntColor <= "000000000000";   -- black
                     
   else 
         cntColor <= "111111111111";   --white background
   end if;
  else
    if((cntHorz < rsec0+35 and cntHorz > lsec0+35 and cntVert < bsec0 and cntVert > tsec0 and value0(charpixcount2)(charpixcount1)='1') 
                       or (cntHorz < rsec1+35 and cntHorz > lsec1+35 and cntVert < bsec1 and cntVert > tsec1 and value1(charpixcount2)(charpixcount1)='1')
                       or (cntHorz < rsec1 and cntHorz > lsec1 and cntVert < bsec1 and cntVert > tsec1 and equal(charpixcount2)(charpixcount1)='1')
                       or (cntHorz < rsec1-35 and cntHorz > lsec1-35 and cntVert < bsec1 and cntVert > tsec1 and ess(charpixcount2)(charpixcount1)='1')
                       or (cntHorz < rsec1-70 and cntHorz > lsec1-70 and cntVert < bsec1 and cntVert > tsec1 and tee(charpixcount2)(charpixcount1)='1')
                       ) then
                       cntColor <= "000000000000";   -- black color for counter display
                       
     else 
           cntColor <= "111111111111";   --white background
     end if;
 
    end if;
    end if;

    end process;

 
     
    vs  <= sncVert;
    hs  <= sncHorz;
    process(blkDisp)
    begin
    if blkDisp ='0' then
    blu <= cntColor(3 downto 0) ;
    grn <= cntColor(7 downto 4) ;
    red <= cntColor(11 downto 8);
    else 
    blu <= "0000";
    grn <= "0000";
    red <= "0000";
    end if;
    end process;
end Behavioral;
